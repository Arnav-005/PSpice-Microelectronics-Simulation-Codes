*Inverting OpAmp
V1 1 0 sin(0 1 1k)
X1 0 2 4 5 3 uA741
R1 1 2 5k
R2 2 3 20K
Vp 4 0 +10V
Vn 5 0 -10V

.lib nom.lib 

.tran 0.01m 4m 0 0.01m
.probe
.end