*RC CIRCUIT
R 2 0 5k
C 1 2 0.1u
V 1 0 AC 1

.AC Dec 20 1 10MEG
.probe
.end