*Astable Multivibrator
X1 2 1 4 5 3 uA741
C1 1 0 0.1u
R1 2 0 10k
R2 2 3 10k
R3 1 3 4.55k
Vp 4 0 +10V
Vn 5 0 -10V

.lib nom.lib

.tran 1u 4m 0 1u
*time period of required square wave is 1m
*stop time of 4m gives 4 cycles

.probe
.end