*Wilson current mirror
V1 6 0 DC 5V
I1 0 5 DC 100mA
R1 5 6 25
Q3 3 2 0 0 npn_transistor_3
Q2 2 2 0 0 npn_transistor_2
Q1 5 3 2 0 npn_transistor_1
.model npn_transistor_1 npn (Is=1.8104e-15 Bf=100) 
.model npn_transistor_2 npn (Is=1.8104e-15 Bf=100) 
.model npn_transistor_3 npn (Is=1.8104e-15 Bf=100) 
.tran 1m 100m 10m�10m
.probe
.end