*RL CIRCUIT
R 1 2 5k
L 2 0 2m
V 1 0 AC 1

.AC Dec 20 1 100MEG
.probe
.end