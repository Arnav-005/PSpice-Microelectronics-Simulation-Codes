*Active HP filter
V1 1 0 AC +1
R1 1 2 10k
C1 2 3 0.01u
R2 3 4 10k
RL 4 0 10k
X1 0 3 5 6 4 uA741
Vp 5 0 +10
Vn 6 0 -10
.lib nom.lib

.ac dec 20 0.01 100k
.probe
.end 