*Difference amplifier
V1 1 0 sin(0 1 1k)
V2 2 0 sin(0 5 1k)
V3 0 6 10
V4 5 0 10

X1 4 3 5 6 7 uA741
R1 3 1 2k
R2 4 2 2k

*attenuating resistors
R3 4 0 4k
R4 7 3 4k

.tran 0.01m 5m 0 0.01m
.lib nom.lib
.probe
.end