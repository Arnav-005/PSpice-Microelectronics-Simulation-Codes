*CE BJT Amplifier
Vsig 1 0 AC 1
Vcc 3 0 +12V
Rb1 2 0 10k
Rb2 2 3 100k
Rc 3 4 20k
Re 5 0 1k
RL 6 0 10k
Cc1 1 2 1u
Cc2 4 6 1u
Ce 5 0 20u
Q1 4 2 5 Q2N2222A
.model Q2N2222A NPN (Is=14.34f Xti=3 Eg=1.11 Vaf=74.03 Bf=255.9 Ne=1.307
+ Ise=14.34f Ikf=.2847 Xtb=1.5 Br=6.092 Nc=2 Isc=0 Ikr=0 Rc=1
+ Cjc=7.306p Mjc=.3416 Vjc=.75 Fc=.5 Cje=22.01p Mje=.377 Vje=.75
+ Tr=46.91n Tf=411.1p Itf=.6 Vtf=1.7 Xtf=3 Rb=10)

.ac oct 10 1 1gig
.probe
.end