*Sallen-key high pass filter 
Vin 1 0 AC 1
R1 3 0 1k
R2 2 4 1k
C2 3 2 0.01u
C1 1 2 0.01u
X1 3 4 5 6 4 UA741
Vp 5 0 DC 10 
Vn 6 0 DC -10
.lib nom.lib 
.ac dec 10 10 500k
.probe 
.end