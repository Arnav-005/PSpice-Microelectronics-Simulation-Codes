*Passive Differentiator
R1 2 0 10k
C1 1 2 0.01u
Vin 1 0 Pulse(0 5 0 0.01f 0.01f 1m 2m)

.tran 0.01m 4m 0 0.01m
.probe
.end