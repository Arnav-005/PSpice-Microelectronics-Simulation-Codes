*MOSFET current mirror
V1 2 0 DC +12
R1 2 1 5
M1 1 1 0 0 nmosfet1
M2 3 1 0 0 nmosfet2
R2 2 3 5

.model nmosfet1 NMOS (LEVEL=3 L=2e-06 W=0.5 KP=2e-05 RS=0.01 
+ RD=0.01 VTO=3 RDS=1000000 TOX=2e-06 CGSO=4e-11 CGDO=1e-11
+ CBD=1e-09 MJ=0.5 PB=0.8 FC=0.5 RG=5 IS=1e-14 N=1 RB=0.001 PHI=0.6
+ GAMMA=0 DELTA=0 ETA=0 THETA=0 KAPPA=0 VMAX=0 XJ=0 UO=600)

.model nmosfet2 NMOS (LEVEL=3 L=2e-06 W=0.5 KP=2e-05 RS=0.01 
+ RD=0.01 VTO=3 RDS=1000000 TOX=2e-06 CGSO=4e-11 CGDO=1e-11
+ CBD=1e-09 MJ=0.5 PB=0.8 FC=0.5 RG=5 IS=1e-14 N=1 RB=0.001 PHI=0.6
+ GAMMA=0 DELTA=0 ETA=0 THETA=0 KAPPA=0 VMAX=0 XJ=0 UO=600)

.tran 0.01m 4m 0 0.01m
.probe
.end