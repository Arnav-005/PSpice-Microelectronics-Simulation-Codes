*OpAmp Freqency Response
X1 1 2 4 5 3 uA741
R1 2 0 10k
R2 2 3 10K
Vp 4 0 +10V
Vn 5 0 -10V
Vin 1 0 AC 1m

.lib nom.lib 

.ac dec 100 1 100meg
.probe
.end